module sin_8bit(input [7:0] bit8_word,
  output reg [7:0] bit8_sin_word);


always @ (*) begin
	case(bit8_word)
		8'b00000000: bit8_sin_word = 8'b10000000;
		8'b00000001: bit8_sin_word = 8'b10000011;
		8'b00000010: bit8_sin_word = 8'b10000110;
		8'b00000011: bit8_sin_word = 8'b10001001;
		8'b00000100: bit8_sin_word = 8'b10001101;
		8'b00000101: bit8_sin_word = 8'b10010000;
		8'b00000110: bit8_sin_word = 8'b10010011;
		8'b00000111: bit8_sin_word = 8'b10010110;
		8'b00001000: bit8_sin_word = 8'b10011001;
		8'b00001001: bit8_sin_word = 8'b10011100;
		8'b00001010: bit8_sin_word = 8'b10011111;
		8'b00001011: bit8_sin_word = 8'b10100010;
		8'b00001100: bit8_sin_word = 8'b10100101;
		8'b00001101: bit8_sin_word = 8'b10101000;
		8'b00001110: bit8_sin_word = 8'b10101011;
		8'b00001111: bit8_sin_word = 8'b10101110;
		8'b00010000: bit8_sin_word = 8'b10110001;
		8'b00010001: bit8_sin_word = 8'b10110100;
		8'b00010010: bit8_sin_word = 8'b10110111;
		8'b00010011: bit8_sin_word = 8'b10111010;
		8'b00010100: bit8_sin_word = 8'b10111100;
		8'b00010101: bit8_sin_word = 8'b10111111;
		8'b00010110: bit8_sin_word = 8'b11000010;
		8'b00010111: bit8_sin_word = 8'b11000100;
		8'b00011000: bit8_sin_word = 8'b11000111;
		8'b00011001: bit8_sin_word = 8'b11001010;
		8'b00011010: bit8_sin_word = 8'b11001100;
		8'b00011011: bit8_sin_word = 8'b11001111;
		8'b00011100: bit8_sin_word = 8'b11010001;
		8'b00011101: bit8_sin_word = 8'b11010100;
		8'b00011110: bit8_sin_word = 8'b11010110;
		8'b00011111: bit8_sin_word = 8'b11011000;
		8'b00100000: bit8_sin_word = 8'b11011011;
		8'b00100001: bit8_sin_word = 8'b11011101;
		8'b00100010: bit8_sin_word = 8'b11011111;
		8'b00100011: bit8_sin_word = 8'b11100001;
		8'b00100100: bit8_sin_word = 8'b11100011;
		8'b00100101: bit8_sin_word = 8'b11100101;
		8'b00100110: bit8_sin_word = 8'b11100111;
		8'b00100111: bit8_sin_word = 8'b11101001;
		8'b00101000: bit8_sin_word = 8'b11101010;
		8'b00101001: bit8_sin_word = 8'b11101100;
		8'b00101010: bit8_sin_word = 8'b11101110;
		8'b00101011: bit8_sin_word = 8'b11101111;
		8'b00101100: bit8_sin_word = 8'b11110001;
		8'b00101101: bit8_sin_word = 8'b11110010;
		8'b00101110: bit8_sin_word = 8'b11110100;
		8'b00101111: bit8_sin_word = 8'b11110101;
		8'b00110000: bit8_sin_word = 8'b11110110;
		8'b00110001: bit8_sin_word = 8'b11110111;
		8'b00110010: bit8_sin_word = 8'b11111001;
		8'b00110011: bit8_sin_word = 8'b11111010;
		8'b00110100: bit8_sin_word = 8'b11111010;
		8'b00110101: bit8_sin_word = 8'b11111011;
		8'b00110110: bit8_sin_word = 8'b11111100;
		8'b00110111: bit8_sin_word = 8'b11111101;
		8'b00111000: bit8_sin_word = 8'b11111110;
		8'b00111001: bit8_sin_word = 8'b11111110;
		8'b00111010: bit8_sin_word = 8'b11111111;
		8'b00111011: bit8_sin_word = 8'b11111111;
		8'b00111100: bit8_sin_word = 8'b11111111;
		8'b00111101: bit8_sin_word = 8'b11111111;
		8'b00111110: bit8_sin_word = 8'b11111111;
		8'b00111111: bit8_sin_word = 8'b11111111;
		8'b01000000: bit8_sin_word = 8'b11111111;
		8'b01000001: bit8_sin_word = 8'b11111111;
		8'b01000010: bit8_sin_word = 8'b11111111;
		8'b01000011: bit8_sin_word = 8'b11111111;
		8'b01000100: bit8_sin_word = 8'b11111111;
		8'b01000101: bit8_sin_word = 8'b11111111;
		8'b01000110: bit8_sin_word = 8'b11111111;
		8'b01000111: bit8_sin_word = 8'b11111110;
		8'b01001000: bit8_sin_word = 8'b11111110;
		8'b01001001: bit8_sin_word = 8'b11111101;
		8'b01001010: bit8_sin_word = 8'b11111100;
		8'b01001011: bit8_sin_word = 8'b11111011;
		8'b01001100: bit8_sin_word = 8'b11111010;
		8'b01001101: bit8_sin_word = 8'b11111010;
		8'b01001110: bit8_sin_word = 8'b11111001;
		8'b01001111: bit8_sin_word = 8'b11110111;
		8'b01010000: bit8_sin_word = 8'b11110110;
		8'b01010001: bit8_sin_word = 8'b11110101;
		8'b01010010: bit8_sin_word = 8'b11110100;
		8'b01010011: bit8_sin_word = 8'b11110010;
		8'b01010100: bit8_sin_word = 8'b11110001;
		8'b01010101: bit8_sin_word = 8'b11101111;
		8'b01010110: bit8_sin_word = 8'b11101110;
		8'b01010111: bit8_sin_word = 8'b11101100;
		8'b01011000: bit8_sin_word = 8'b11101010;
		8'b01011001: bit8_sin_word = 8'b11101001;
		8'b01011010: bit8_sin_word = 8'b11100111;
		8'b01011011: bit8_sin_word = 8'b11100101;
		8'b01011100: bit8_sin_word = 8'b11100011;
		8'b01011101: bit8_sin_word = 8'b11100001;
		8'b01011110: bit8_sin_word = 8'b11011111;
		8'b01011111: bit8_sin_word = 8'b11011101;
		8'b01100000: bit8_sin_word = 8'b11011011;
		8'b01100001: bit8_sin_word = 8'b11011000;
		8'b01100010: bit8_sin_word = 8'b11010110;
		8'b01100011: bit8_sin_word = 8'b11010100;
		8'b01100100: bit8_sin_word = 8'b11010001;
		8'b01100101: bit8_sin_word = 8'b11001111;
		8'b01100110: bit8_sin_word = 8'b11001100;
		8'b01100111: bit8_sin_word = 8'b11001010;
		8'b01101000: bit8_sin_word = 8'b11000111;
		8'b01101001: bit8_sin_word = 8'b11000100;
		8'b01101010: bit8_sin_word = 8'b11000010;
		8'b01101011: bit8_sin_word = 8'b10111111;
		8'b01101100: bit8_sin_word = 8'b10111100;
		8'b01101101: bit8_sin_word = 8'b10111010;
		8'b01101110: bit8_sin_word = 8'b10110111;
		8'b01101111: bit8_sin_word = 8'b10110100;
		8'b01110000: bit8_sin_word = 8'b10110001;
		8'b01110001: bit8_sin_word = 8'b10101110;
		8'b01110010: bit8_sin_word = 8'b10101011;
		8'b01110011: bit8_sin_word = 8'b10101000;
		8'b01110100: bit8_sin_word = 8'b10100101;
		8'b01110101: bit8_sin_word = 8'b10100010;
		8'b01110110: bit8_sin_word = 8'b10011111;
		8'b01110111: bit8_sin_word = 8'b10011100;
		8'b01111000: bit8_sin_word = 8'b10011001;
		8'b01111001: bit8_sin_word = 8'b10010110;
		8'b01111010: bit8_sin_word = 8'b10010011;
		8'b01111011: bit8_sin_word = 8'b10010000;
		8'b01111100: bit8_sin_word = 8'b10001101;
		8'b01111101: bit8_sin_word = 8'b10001001;
		8'b01111110: bit8_sin_word = 8'b10000110;
		8'b01111111: bit8_sin_word = 8'b10000011;
		8'b10000000: bit8_sin_word = 8'b10000000;
		8'b10000001: bit8_sin_word = 8'b01111101;
		8'b10000010: bit8_sin_word = 8'b01111010;
		8'b10000011: bit8_sin_word = 8'b01110111;
		8'b10000100: bit8_sin_word = 8'b01110011;
		8'b10000101: bit8_sin_word = 8'b01110000;
		8'b10000110: bit8_sin_word = 8'b01101101;
		8'b10000111: bit8_sin_word = 8'b01101010;
		8'b10001000: bit8_sin_word = 8'b01100111;
		8'b10001001: bit8_sin_word = 8'b01100100;
		8'b10001010: bit8_sin_word = 8'b01100001;
		8'b10001011: bit8_sin_word = 8'b01011110;
		8'b10001100: bit8_sin_word = 8'b01011011;
		8'b10001101: bit8_sin_word = 8'b01011000;
		8'b10001110: bit8_sin_word = 8'b01010101;
		8'b10001111: bit8_sin_word = 8'b01010010;
		8'b10010000: bit8_sin_word = 8'b01001111;
		8'b10010001: bit8_sin_word = 8'b01001100;
		8'b10010010: bit8_sin_word = 8'b01001001;
		8'b10010011: bit8_sin_word = 8'b01000110;
		8'b10010100: bit8_sin_word = 8'b01000100;
		8'b10010101: bit8_sin_word = 8'b01000001;
		8'b10010110: bit8_sin_word = 8'b00111110;
		8'b10010111: bit8_sin_word = 8'b00111100;
		8'b10011000: bit8_sin_word = 8'b00111001;
		8'b10011001: bit8_sin_word = 8'b00110110;
		8'b10011010: bit8_sin_word = 8'b00110100;
		8'b10011011: bit8_sin_word = 8'b00110001;
		8'b10011100: bit8_sin_word = 8'b00101111;
		8'b10011101: bit8_sin_word = 8'b00101100;
		8'b10011110: bit8_sin_word = 8'b00101010;
		8'b10011111: bit8_sin_word = 8'b00101000;
		8'b10100000: bit8_sin_word = 8'b00100101;
		8'b10100001: bit8_sin_word = 8'b00100011;
		8'b10100010: bit8_sin_word = 8'b00100001;
		8'b10100011: bit8_sin_word = 8'b00011111;
		8'b10100100: bit8_sin_word = 8'b00011101;
		8'b10100101: bit8_sin_word = 8'b00011011;
		8'b10100110: bit8_sin_word = 8'b00011001;
		8'b10100111: bit8_sin_word = 8'b00010111;
		8'b10101000: bit8_sin_word = 8'b00010110;
		8'b10101001: bit8_sin_word = 8'b00010100;
		8'b10101010: bit8_sin_word = 8'b00010010;
		8'b10101011: bit8_sin_word = 8'b00010001;
		8'b10101100: bit8_sin_word = 8'b00001111;
		8'b10101101: bit8_sin_word = 8'b00001110;
		8'b10101110: bit8_sin_word = 8'b00001100;
		8'b10101111: bit8_sin_word = 8'b00001011;
		8'b10110000: bit8_sin_word = 8'b00001010;
		8'b10110001: bit8_sin_word = 8'b00001001;
		8'b10110010: bit8_sin_word = 8'b00000111;
		8'b10110011: bit8_sin_word = 8'b00000110;
		8'b10110100: bit8_sin_word = 8'b00000110;
		8'b10110101: bit8_sin_word = 8'b00000101;
		8'b10110110: bit8_sin_word = 8'b00000100;
		8'b10110111: bit8_sin_word = 8'b00000011;
		8'b10111000: bit8_sin_word = 8'b00000010;
		8'b10111001: bit8_sin_word = 8'b00000010;
		8'b10111010: bit8_sin_word = 8'b00000001;
		8'b10111011: bit8_sin_word = 8'b00000001;
		8'b10111100: bit8_sin_word = 8'b00000001;
		8'b10111101: bit8_sin_word = 8'b00000000;
		8'b10111110: bit8_sin_word = 8'b00000000;
		8'b10111111: bit8_sin_word = 8'b00000000;
		8'b11000000: bit8_sin_word = 8'b00000000;
		8'b11000001: bit8_sin_word = 8'b00000000;
		8'b11000010: bit8_sin_word = 8'b00000000;
		8'b11000011: bit8_sin_word = 8'b00000000;
		8'b11000100: bit8_sin_word = 8'b00000001;
		8'b11000101: bit8_sin_word = 8'b00000001;
		8'b11000110: bit8_sin_word = 8'b00000001;
		8'b11000111: bit8_sin_word = 8'b00000010;
		8'b11001000: bit8_sin_word = 8'b00000010;
		8'b11001001: bit8_sin_word = 8'b00000011;
		8'b11001010: bit8_sin_word = 8'b00000100;
		8'b11001011: bit8_sin_word = 8'b00000101;
		8'b11001100: bit8_sin_word = 8'b00000110;
		8'b11001101: bit8_sin_word = 8'b00000110;
		8'b11001110: bit8_sin_word = 8'b00000111;
		8'b11001111: bit8_sin_word = 8'b00001001;
		8'b11010000: bit8_sin_word = 8'b00001010;
		8'b11010001: bit8_sin_word = 8'b00001011;
		8'b11010010: bit8_sin_word = 8'b00001100;
		8'b11010011: bit8_sin_word = 8'b00001110;
		8'b11010100: bit8_sin_word = 8'b00001111;
		8'b11010101: bit8_sin_word = 8'b00010001;
		8'b11010110: bit8_sin_word = 8'b00010010;
		8'b11010111: bit8_sin_word = 8'b00010100;
		8'b11011000: bit8_sin_word = 8'b00010110;
		8'b11011001: bit8_sin_word = 8'b00010111;
		8'b11011010: bit8_sin_word = 8'b00011001;
		8'b11011011: bit8_sin_word = 8'b00011011;
		8'b11011100: bit8_sin_word = 8'b00011101;
		8'b11011101: bit8_sin_word = 8'b00011111;
		8'b11011110: bit8_sin_word = 8'b00100001;
		8'b11011111: bit8_sin_word = 8'b00100011;
		8'b11100000: bit8_sin_word = 8'b00100101;
		8'b11100001: bit8_sin_word = 8'b00101000;
		8'b11100010: bit8_sin_word = 8'b00101010;
		8'b11100011: bit8_sin_word = 8'b00101100;
		8'b11100100: bit8_sin_word = 8'b00101111;
		8'b11100101: bit8_sin_word = 8'b00110001;
		8'b11100110: bit8_sin_word = 8'b00110100;
		8'b11100111: bit8_sin_word = 8'b00110110;
		8'b11101000: bit8_sin_word = 8'b00111001;
		8'b11101001: bit8_sin_word = 8'b00111100;
		8'b11101010: bit8_sin_word = 8'b00111110;
		8'b11101011: bit8_sin_word = 8'b01000001;
		8'b11101100: bit8_sin_word = 8'b01000100;
		8'b11101101: bit8_sin_word = 8'b01000110;
		8'b11101110: bit8_sin_word = 8'b01001001;
		8'b11101111: bit8_sin_word = 8'b01001100;
		8'b11110000: bit8_sin_word = 8'b01001111;
		8'b11110001: bit8_sin_word = 8'b01010010;
		8'b11110010: bit8_sin_word = 8'b01010101;
		8'b11110011: bit8_sin_word = 8'b01011000;
		8'b11110100: bit8_sin_word = 8'b01011011;
		8'b11110101: bit8_sin_word = 8'b01011110;
		8'b11110110: bit8_sin_word = 8'b01100001;
		8'b11110111: bit8_sin_word = 8'b01100100;
		8'b11111000: bit8_sin_word = 8'b01100111;
		8'b11111001: bit8_sin_word = 8'b01101010;
		8'b11111010: bit8_sin_word = 8'b01101101;
		8'b11111011: bit8_sin_word = 8'b01110000;
		8'b11111100: bit8_sin_word = 8'b01110011;
		8'b11111101: bit8_sin_word = 8'b01110111;
		8'b11111110: bit8_sin_word = 8'b01111010;
		8'b11111111: bit8_sin_word = 8'b01111101;
	endcase
	end
endmodule

